module addition_stage4#
(
    parameter integer 
)
(
    input
    
);

endmodule