`timescale 1ns / 1ps



module fpu_division(
    input [31:0] float_num1,
    input [31:0] float_num2,
    output reg [31:0] div_result,
    output [7:0]pos,
    output sign_out,
    output [47:0] div_out
);

// Partition of floating-point numbers
wire [7:0] exp_num1, exp_num2;
wire [23:0] mantissa_num1, mantissa_num2;
wire sign_num1, sign_num2;

// Outputs from various components
wire [8:0] exponent_subtract;
wire [7:0] adjusted_exponent;

// Normalizer outputs
reg [7:0] normalized_exponent; // Initialize to avoid unset bits
reg [22:0] normalized_mantissa;   // Initialize to avoid unset bits

// Assign input partitions 
assign sign_num1 = float_num1[31];
assign exp_num1 = float_num1[30:23];
assign sign_num2 = float_num2[31];
assign exp_num2 = float_num2[30:23];

// Ensure mantissa is set correctly
assign mantissa_num1 =  {1'b1, float_num1[22:0]};
assign mantissa_num2 =  {1'b1, float_num2[22:0]};

// Exponent difference calculation
assign exponent_subtract = exp_num1 - exp_num2;  // Direct subtraction

// Adjust the exponent (bias correction of 127)
assign adjusted_exponent = exponent_subtract + 8'b0111_1111 ;  // Keep only 8 bits

// Mantissa division result (48-bit precision)
wire [23:0] mantissa_div_result;  
reg [5:0] position;  // 8-bit position
reg [47:0] shifted_mantissa;  
  

nph_divider d0(.mantissa_num1(mantissa_num1),.mantissa_num2(mantissa_num2),.mantissa_div_result(mantissa_div_result));
//assign mantissa_div_result = mantissa_num1 / mantissa_num2;
assign div_out = mantissa_div_result;

always @(*) begin
   
    casez(mantissa_div_result)
        48'b1??????????????????????????????????????????????? : position = 6'd0;
        48'b01?????????????????????????????????????????????? : position = 6'd1;
        48'b001????????????????????????????????????????????? : position = 6'd2;
        48'b0001???????????????????????????????????????????? : position = 6'd3;
        48'b00001??????????????????????????????????????????? : position = 6'd4;
        48'b000001?????????????????????????????????????????? : position = 6'd5;
        48'b0000001????????????????????????????????????????? : position = 6'd6;
        48'b00000001???????????????????????????????????????? : position = 6'd7;
        48'b000000001??????????????????????????????????????? : position = 6'd8;
        48'b0000000001?????????????????????????????????????? : position = 6'd9;
        48'b00000000001????????????????????????????????????? : position = 6'd10;
        48'b000000000001???????????????????????????????????? : position = 6'd11;
        48'b0000000000001??????????????????????????????????? : position = 6'd12;
        48'b00000000000001?????????????????????????????????? : position = 6'd13;
        48'b000000000000001????????????????????????????????? : position = 6'd14;
        48'b0000000000000001???????????????????????????????? : position = 6'd15;
        48'b00000000000000001??????????????????????????????? : position = 6'd16;
        48'b000000000000000001?????????????????????????????? : position = 6'd17;
        48'b0000000000000000001????????????????????????????? : position = 6'd18;
        48'b00000000000000000001???????????????????????????? : position = 6'd19;
        48'b000000000000000000001??????????????????????????? : position = 6'd20;
        48'b0000000000000000000001?????????????????????????? : position = 6'd21;
        48'b00000000000000000000001????????????????????????? : position = 6'd22;
        48'b000000000000000000000001???????????????????????? : position = 6'd23;
        48'b0000000000000000000000001??????????????????????? : position = 6'd24;
        48'b00000000000000000000000001?????????????????????? : position = 6'd25;
        48'b000000000000000000000000001????????????????????? : position = 6'd26;
        48'b0000000000000000000000000001???????????????????? : position = 6'd27;
        48'b00000000000000000000000000001??????????????????? : position = 6'd28;
        48'b000000000000000000000000000001?????????????????? : position = 6'd29;
        48'b0000000000000000000000000000001????????????????? : position = 6'd30;
        48'b00000000000000000000000000000001???????????????? : position = 6'd31;
        48'b000000000000000000000000000000001??????????????? : position = 6'd32;
        48'b0000000000000000000000000000000001?????????????? : position = 6'd33;
        48'b00000000000000000000000000000000001????????????? : position = 6'd34;
        48'b000000000000000000000000000000000001???????????? : position = 6'd35;
        48'b0000000000000000000000000000000000001??????????? : position = 6'd36;
        48'b00000000000000000000000000000000000001?????????? : position = 6'd37;
        48'b000000000000000000000000000000000000001????????? : position = 6'd38;
        48'b0000000000000000000000000000000000000001???????? : position = 6'd39;
        48'b00000000000000000000000000000000000000001??????? : position = 6'd40;
        48'b000000000000000000000000000000000000000001?????? : position = 6'd41;
        48'b0000000000000000000000000000000000000000001????? : position = 6'd42;
        48'b00000000000000000000000000000000000000000001???? : position = 6'd43;
        48'b000000000000000000000000000000000000000000001??? : position = 6'd44;
        48'b0000000000000000000000000000000000000000000001?? : position = 6'd45;
        48'b00000000000000000000000000000000000000000000001? : position = 6'd46;
        48'b000000000000000000000000000000000000000000000001 : position = 6'd47;
        default: position = 6'd48; // No bits set, assume denormalized
    endcase
end

//// Normalize Mantissa and Exponent
always @(*) begin
   
        shifted_mantissa = mantissa_div_result << position;  
        normalized_mantissa = shifted_mantissa[47:25];  // Take upper 23 bits
        normalized_exponent = adjusted_exponent;  
end

assign pos = position;

// Calculate the output sign

assign  sign_out = float_num1[31] ^float_num2[31];


// Combine the final result
always @(*) begin
    div_result = {sign_out, normalized_exponent, normalized_mantissa};
end

endmodule
