`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/02/2025 12:37:04 PM
// Design Name: 
// Module Name: mutliplication
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mutliplication
#(parameter D_WIDTH = 32,
  parameter M_WIDTH = 23,
  parameter E_WIDTH = 8
 )
 (
    input  [D_WIDTH-1 : 0]number_1,
    input  [D_WIDTH-1 : 0]number_2,
    output [D_WIDTH-1 : 0]number_out,
    output [E_WIDTH-1:0]pos  
 );
    //Partitioning bits for sign,exponent,mantissa;
    wire                sign1,sign2;
    wire [E_WIDTH-1 : 0]exp1,exp2;
    wire [M_WIDTH-1 : 0]m1,m2;
    
    //Final sign, exponent and mantissa
    wire [E_WIDTH-1 : 0]output_exponent;
    wire [M_WIDTH-1 : 0]output_mantissa;
    wire                output_sign;
    
    //input Numbers
    assign sign1 = number_1[D_WIDTH-1]; //[31]
    assign exp1  = number_1[D_WIDTH-2 -: E_WIDTH]; //[30:23]
    assign m1    = number_1[M_WIDTH-1 -: M_WIDTH]; //[22:0]
    
    assign sign2 = number_2[D_WIDTH-1];
    assign exp2  = number_2[D_WIDTH-2 -: E_WIDTH];
    assign m2    = number_2[M_WIDTH-1 -: M_WIDTH];
    
    //Intermediate outputs
    wire [E_WIDTH : 0]exp_out;
    wire [E_WIDTH : 0]unbiased_exp_out;
    wire [47:0]multiply_out;
    
    //Input for passing to the normalizer
    reg [47:0]mantissa;
    reg [47:0]shifted_mantissa;
    
    reg [7:0]position;
    
    //Outputs from the normalizer
    reg [47:0]normalized_mantissa;
    reg [8:0] normalized_exponent;
    
    // Exponent Addition
    assign exp_out = exp1 + exp2;
    
    //Unbiasing the exp_out with 127
    assign unbiased_exp_out = exp_out - 8'b0111_1111;
    
    //Multiplying the mantissas
    assign multiply_out = {1'b1, m1} * {1'b1 ,m2};
    
    //Normalizer_Part
    always @ (*)
    begin
        mantissa = multiply_out;
        
        casez(mantissa)
        48'b1??????????????????????????????????????????????? : position = 8'd0;
        48'b01?????????????????????????????????????????????? : position = 8'd1;
        48'b001????????????????????????????????????????????? : position = 8'd2;
        48'b0001???????????????????????????????????????????? : position = 8'd3;
        48'b00001??????????????????????????????????????????? : position = 8'd4;
        48'b000001?????????????????????????????????????????? : position = 8'd5;
        48'b0000001????????????????????????????????????????? : position = 8'd6;
        48'b00000001???????????????????????????????????????? : position = 8'd7;
        48'b000000001??????????????????????????????????????? : position = 8'd8;
        48'b0000000001?????????????????????????????????????? : position = 8'd9;
        48'b00000000001????????????????????????????????????? : position = 8'd10;
        48'b000000000001???????????????????????????????????? : position = 8'd11;
        48'b0000000000001??????????????????????????????????? : position = 8'd12;
        48'b00000000000001?????????????????????????????????? : position = 8'd13;
        48'b000000000000001????????????????????????????????? : position = 8'd14;
        48'b0000000000000001???????????????????????????????? : position = 8'd15;
        48'b00000000000000001??????????????????????????????? : position = 8'd16;
        48'b000000000000000001?????????????????????????????? : position = 8'd17;
        48'b0000000000000000001????????????????????????????? : position = 8'd18;
        48'b00000000000000000001???????????????????????????? : position = 8'd19;
        48'b000000000000000000001??????????????????????????? : position = 8'd20;
        48'b0000000000000000000001?????????????????????????? : position = 8'd21;
        48'b00000000000000000000001????????????????????????? : position = 8'd22;
        48'b000000000000000000000001???????????????????????? : position = 8'd23;
        default: position = 8'd24; // Assume denormalized
        endcase
    end
    assign pos = position;
    
    //Mantissa Alignment for final output
    always @ (*)
    begin
        shifted_mantissa = mantissa << (position + 1);
        normalized_mantissa = shifted_mantissa[47:25];
        normalized_exponent = (unbiased_exp_out - position) + 1;
    end
    
    assign output_mantissa = normalized_mantissa;
    assign output_exponent = normalized_exponent;
    assign output_sign     = sign1 ^ sign2;
    
    //Final Result
    assign number_out = {output_sign, output_exponent, output_mantissa};
    
endmodule
