module floating_point_addition#
(
    parameter integer DATA_WIDTH = 32
)
(
    input  [DATA_WIDTH-1:0] floating1,
    input  [DATA_WIDTH-1:0] floating2,

    output [DATA_WIDTH-1:0] floating_addition_out
);

    wire sign1,sign2;
    wire [DATA_WIDTH-1:0]mentissa1,mentissa2;
    
endmodule